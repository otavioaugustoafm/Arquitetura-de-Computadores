/*Guia_0201.v851568 - Otávio Augusto de Assis Ferreira Monteiro*/module Guia_020a;// define datareal x = 0 ; // decimalreal power2 = 1.0; // power of 2integer y = 4 ; // counterreg [4:0] b = 5'b00011; // binary (only fraction part, Big Endian)// actionsinitialbegin : main$display ( "Guia_0201 - Tests" );while ( y >= 0 )beginpower2 = power2 / 2.0;if ( b[y] == 1 )beginx = x + power2;endy=y-1;end // end whilex = x + 0;$display ( "a) = %f", x);end // mainendmodule // Guia_0201amodule Guia_020b;// define datareal x = 0 ; // decimalreal power2 = 1.0; // power of 2integer y = 4 ; // counterreg [4:0] b = 5'b01001; // binary (only fraction part, Big Endian)// actionsinitialbegin : mainwhile ( y >= 0 )beginpower2 = power2 / 2.0;if ( b[y] == 1 )beginx = x + power2;endy=y-1;end // end whilex = x + 0;$display ( "b) = %f", x);end // mainendmodule // Guia_0201bmodule Guia_020c;// define datareal x = 0 ; // decimalreal power2 = 1.0; // power of 2integer y = 4 ; // counterreg [4:0] b = 5'b10101; // binary (only fraction part, Big Endian)// actionsinitialbegin : mainwhile ( y >= 0 )beginpower2 = power2 / 2.0;if ( b[y] == 1 )beginx = x + power2;endy=y-1;end // end whilex = x + 0;$display ( "c) = %f", x);end // mainendmodule // Guia_0201cmodule Guia_020d;// define datareal x = 0 ; // decimalreal power2 = 1.0; // power of 2integer y = 4 ; // counterreg [4:0] b = 5'b11101; // binary (only fraction part, Big Endian)// actionsinitialbegin : mainwhile ( y >= 0 )beginpower2 = power2 / 2.0;if ( b[y] == 1 )beginx = x + power2;endy=y-1;end // end whilex = x + 1;$display ( "d) = %f", x);end // mainendmodule // Guia_0201dmodule Guia_020e;// define datareal x = 0 ; // decimalreal power2 = 1.0; // power of 2integer y = 4 ; // counterreg [4:0] b = 5'b11001; // binary (only fraction part, Big Endian)// actionsinitialbegin : mainwhile ( y >= 0 )beginpower2 = power2 / 2.0;if ( b[y] == 1 )beginx = x + power2;endy=y-1;end // end whilex = x + 3;$display ( "e) = %f", x);end // mainendmodule // Guia_0201e